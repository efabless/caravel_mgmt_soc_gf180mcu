VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180_ram_512x8_wrapper
  CLASS BLOCK ;
  FOREIGN gf180_ram_512x8_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 444.860 BY 512.880 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 508.880 252.560 512.880 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 508.880 259.280 512.880 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 508.880 266.000 512.880 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 508.880 158.480 512.880 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 508.880 165.200 512.880 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 508.880 171.920 512.880 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 508.880 178.640 512.880 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 508.880 272.720 512.880 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 508.880 279.440 512.880 ;
    END
  END A[8]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 508.880 185.360 512.880 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 508.880 286.160 512.880 ;
    END
  END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 508.880 420.560 512.880 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 508.880 380.240 512.880 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 508.880 360.080 512.880 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 508.880 306.320 512.880 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 508.880 138.320 512.880 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 508.880 84.560 512.880 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 508.880 64.400 512.880 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 508.880 17.360 512.880 ;
    END
  END D[7]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 508.880 225.680 512.880 ;
    END
  END GWEN
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 508.880 407.120 512.880 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 508.880 386.960 512.880 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 508.880 353.360 512.880 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 508.880 319.760 512.880 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 508.880 124.880 512.880 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 508.880 91.280 512.880 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 508.880 57.680 512.880 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 508.880 30.800 512.880 ;
    END
  END Q[7]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 5.220 15.680 8.220 493.920 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 428.630 15.680 431.630 493.920 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.22 14.18 437.92 17.18 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 9.220 15.680 12.220 493.920 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 432.630 15.680 435.630 493.920 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.72 18.18 437.92 21.18 ;
    END
  END VSS
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 508.880 413.840 512.880 ;
    END
  END WEN[0]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 508.880 373.520 512.880 ;
    END
  END WEN[1]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 508.880 366.800 512.880 ;
    END
  END WEN[2]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 508.880 313.040 512.880 ;
    END
  END WEN[3]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 508.880 131.600 512.880 ;
    END
  END WEN[4]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 508.880 77.840 512.880 ;
    END
  END WEN[5]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 508.880 71.120 512.880 ;
    END
  END WEN[6]
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 508.880 24.080 512.880 ;
    END
  END WEN[7]
  OBS
      LAYER Metal1 ;
        RECT 5.000 5.000 436.860 489.880 ;
      LAYER Metal2 ;
        RECT 5.000 508.580 16.500 509.460 ;
        RECT 17.660 508.580 23.220 509.460 ;
        RECT 24.380 508.580 29.940 509.460 ;
        RECT 31.100 508.580 56.820 509.460 ;
        RECT 57.980 508.580 63.540 509.460 ;
        RECT 64.700 508.580 70.260 509.460 ;
        RECT 71.420 508.580 76.980 509.460 ;
        RECT 78.140 508.580 83.700 509.460 ;
        RECT 84.860 508.580 90.420 509.460 ;
        RECT 91.580 508.580 124.020 509.460 ;
        RECT 125.180 508.580 130.740 509.460 ;
        RECT 131.900 508.580 137.460 509.460 ;
        RECT 138.620 508.580 157.620 509.460 ;
        RECT 158.780 508.580 164.340 509.460 ;
        RECT 165.500 508.580 171.060 509.460 ;
        RECT 172.220 508.580 177.780 509.460 ;
        RECT 178.940 508.580 184.500 509.460 ;
        RECT 185.660 508.580 224.820 509.460 ;
        RECT 225.980 508.580 251.700 509.460 ;
        RECT 252.860 508.580 258.420 509.460 ;
        RECT 259.580 508.580 265.140 509.460 ;
        RECT 266.300 508.580 271.860 509.460 ;
        RECT 273.020 508.580 278.580 509.460 ;
        RECT 279.740 508.580 285.300 509.460 ;
        RECT 286.460 508.580 305.460 509.460 ;
        RECT 306.620 508.580 312.180 509.460 ;
        RECT 313.340 508.580 318.900 509.460 ;
        RECT 320.060 508.580 352.500 509.460 ;
        RECT 353.660 508.580 359.220 509.460 ;
        RECT 360.380 508.580 365.940 509.460 ;
        RECT 367.100 508.580 372.660 509.460 ;
        RECT 373.820 508.580 379.380 509.460 ;
        RECT 380.540 508.580 386.100 509.460 ;
        RECT 387.260 508.580 406.260 509.460 ;
        RECT 407.420 508.580 412.980 509.460 ;
        RECT 414.140 508.580 419.700 509.460 ;
        RECT 420.860 508.580 436.860 509.460 ;
        RECT 5.000 5.000 436.860 508.580 ;
      LAYER Metal3 ;
        RECT 5.000 5.000 436.860 504.980 ;
  END
END gf180_ram_512x8_wrapper
END LIBRARY

