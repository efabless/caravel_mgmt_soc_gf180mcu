VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180_ram_512x8_wrapper
  CLASS BLOCK ;
  FOREIGN gf180_ram_512x8_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 444.860 BY 495.880 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.720 491.880 265.280 495.880 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.220 491.880 273.780 495.880 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.720 491.880 282.280 495.880 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.720 491.880 155.280 495.880 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.720 491.880 160.280 495.880 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.720 491.880 164.280 495.880 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.720 491.880 167.280 495.880 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.220 491.880 287.780 495.880 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.720 491.880 291.280 495.880 ;
    END
  END A[8]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.220 491.880 184.780 495.880 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.220 491.880 296.780 495.880 ;
    END
  END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 491.880 427.280 495.880 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.720 491.880 375.280 495.880 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 368.720 491.880 369.280 495.880 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.720 491.880 317.280 495.880 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.720 491.880 129.280 495.880 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.220 491.880 77.780 495.880 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.720 491.880 71.280 495.880 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 18.720 491.880 19.280 495.880 ;
    END
  END D[7]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.840 491.880 233.400 495.880 ;
    END
  END GWEN
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 419.220 491.880 419.780 495.880 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.220 491.880 378.780 495.880 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.220 491.880 365.780 495.880 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.720 491.880 325.280 495.880 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.220 491.880 121.780 495.880 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.220 491.880 80.780 495.880 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.220 491.880 67.780 495.880 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.720 491.880 27.280 495.880 ;
    END
  END Q[7]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 5.220 14.180 8.220 478.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 428.630 14.180 431.630 478.240 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.220 14.180 437.920 17.180 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 9.220 15.680 12.220 478.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 432.630 15.680 435.630 478.240 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.720 18.180 437.920 21.180 ;
    END
  END VSS
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.220 491.880 423.780 495.880 ;
    END
  END WEN[0]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.720 491.880 373.280 495.880 ;
    END
  END WEN[1]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 491.880 371.280 495.880 ;
    END
  END WEN[2]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.720 491.880 319.280 495.880 ;
    END
  END WEN[3]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 125.220 491.880 125.780 495.880 ;
    END
  END WEN[4]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 74.970 491.880 75.530 495.880 ;
    END
  END WEN[5]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.720 491.880 73.280 495.880 ;
    END
  END WEN[6]
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.220 491.880 22.780 495.880 ;
    END
  END WEN[7]
  OBS
      LAYER Metal1 ;
        RECT 5.000 5.000 436.860 489.880 ;
      LAYER Metal2 ;
        RECT 5.000 491.580 18.420 492.520 ;
        RECT 19.580 491.580 21.920 492.520 ;
        RECT 23.080 491.580 26.420 492.520 ;
        RECT 27.580 491.580 66.920 492.520 ;
        RECT 68.080 491.580 70.420 492.520 ;
        RECT 71.580 491.580 72.420 492.520 ;
        RECT 73.580 491.580 74.670 492.520 ;
        RECT 75.830 491.580 76.920 492.520 ;
        RECT 78.080 491.580 79.920 492.520 ;
        RECT 81.080 491.580 120.920 492.520 ;
        RECT 122.080 491.580 124.920 492.520 ;
        RECT 126.080 491.580 128.420 492.520 ;
        RECT 129.580 491.580 154.420 492.520 ;
        RECT 155.580 491.580 159.420 492.520 ;
        RECT 160.580 491.580 163.420 492.520 ;
        RECT 164.580 491.580 166.420 492.520 ;
        RECT 167.580 491.580 183.920 492.520 ;
        RECT 185.080 491.580 232.540 492.520 ;
        RECT 233.700 491.580 264.420 492.520 ;
        RECT 265.580 491.580 272.920 492.520 ;
        RECT 274.080 491.580 281.420 492.520 ;
        RECT 282.580 491.580 286.920 492.520 ;
        RECT 288.080 491.580 290.420 492.520 ;
        RECT 291.580 491.580 295.920 492.520 ;
        RECT 297.080 491.580 316.420 492.520 ;
        RECT 317.580 491.580 318.420 492.520 ;
        RECT 319.580 491.580 324.420 492.520 ;
        RECT 325.580 491.580 364.920 492.520 ;
        RECT 366.080 491.580 368.420 492.520 ;
        RECT 369.580 491.580 370.420 492.520 ;
        RECT 371.580 491.580 372.420 492.520 ;
        RECT 373.580 491.580 374.420 492.520 ;
        RECT 375.580 491.580 377.920 492.520 ;
        RECT 379.080 491.580 418.920 492.520 ;
        RECT 420.080 491.580 422.920 492.520 ;
        RECT 424.080 491.580 426.420 492.520 ;
        RECT 427.580 491.580 436.860 492.520 ;
        RECT 5.000 5.000 436.860 491.580 ;
      LAYER Metal3 ;
        RECT 5.000 5.000 436.860 489.880 ;
  END
END gf180_ram_512x8_wrapper
END LIBRARY

